module gray2bin
  #(parameter width_p = 5)
   // You must fill these in with width_p
   (input [width_p-1:0] gray_i
    ,output [width_p-1:0] bin_o);

  logic [width_p-1:0] bin_l;

  always_comb begin
    bin_l[width_p-1] = gray_i[width_p-1];
    for (int i = width_p-2; i >= 0; i--) begin
      bin_l[i] = bin_l[i+1] ^ gray_i[i];
    end
  end
  
  assign bin_o = bin_l;

endmodule
