module full_add
  (input [0:0] a_i
  ,input [0:0] b_i
  ,input [0:0] carry_i
  ,output [0:0] carry_o
  ,output [0:0] sum_o);

   // For Lab 2, you may use assign statements!
   // Your code here:

  logic [0:0] sum_l;
  logic [0:0] carry_l;

  always_comb begin
    sum_l = a_i ^ b_i ^ carry_i;
    carry_l = (a_i & b_i) | (b_i & carry_i) | (a_i & carry_i);
  end

  assign sum_o = sum_l;
  assign carry_o = carry_l;

endmodule
